** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/VCO_tb.sch
**.subckt VCO_tb
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
XM1 VBIAS VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM2 VBIAS VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
V4 net1 VSS 2
.save i(v4)
C2 VBIAS VSS 1p m=1
V3 VCTRL VSS pwl(0 0 0.1n 1 100n 1 101n 2 120n 2 121n 3)
.save i(v3)
xVCO1 VDD VSS VBIAS VCTRL net3 VCO
xinv_one1 VDD VSS net3 net2 INV_one
xinv_four1 VDD VSS net2 OUT INV_four
C1 OUT VSS 10f m=1
**** begin user architecture code

.include /home/shahidosic/OSPDKs/GF180/PDK/share/pdk/gf180mcuC/libs.tech/ngspice/design.spice
.lib /home/shahidosic/OSPDKs/GF180/PDK/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.spice typical



.ic v(OUT)=0
.option TEMP=27
.control
save all
tran 10p 150n
plot v(VCTRL) v(OUT)
write inv_tb.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/VCO.sym # of pins=5
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/VCO.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/VCO.sch
.subckt VCO VDD VSS VBIAS VCTRL OSC
*.iopin VDD
*.iopin VSS
*.iopin OSC
*.iopin VBIAS
*.iopin VCTRL
XM5 net7 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM3 net8 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM4 net9 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM8 net10 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM9 net11 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM10 net12 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM11 net13 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM6 net14 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM7 net15 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM12 net16 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM13 net17 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM15 net18 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM16 net19 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM17 net20 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
xinv1 net7 net14 OSC net1 inv
xinv2 net8 net15 net1 net2 inv
xinv3 net9 net16 net2 net3 inv
xinv4 net10 net17 net3 net4 inv
xinv5 net11 net18 net4 net5 inv
xinv6 net12 net19 net5 net6 inv
xinv7 net13 net20 net6 OSC inv
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/INV_one.sym # of pins=4
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/INV_one.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/INV_one.sch
.subckt INV_one VDD VSS IN OUT
*.ipin IN
*.iopin VDD
*.iopin VSS
*.opin OUT
XM1 OUT IN VSS VSS nmos_3p3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/INV_four.sym # of pins=4
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/INV_four.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/INV_four.sch
.subckt INV_four VDD VSS IN OUT
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
xinv_one1 VDD VSS IN OUT INV_one
xinv_one2 VDD VSS IN OUT INV_one
xinv_one3 VDD VSS IN OUT INV_one
xinv_one4 VDD VSS IN OUT INV_one
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/inv.sym # of pins=4
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/inv.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/inv.sch
.subckt inv VDD VSS IN OUT
*.ipin IN
*.iopin VDD
*.iopin VSS
*.opin OUT
XM1 OUT IN VSS VSS nmos_3p3 L=1u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM2 OUT IN VDD VDD pmos_3p3 L=1u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
.ends

.GLOBAL GND
.end
