** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/Oscillator.sch
**.subckt Oscillator
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3
.save i(v2)
xTest_INV1 VDD VSS OUT net1 Test_INV
xTest_INV2 VDD VSS net1 net2 Test_INV
xTest_INV3 VDD VSS net2 net3 Test_INV
xTest_INV4 VDD VSS net3 net4 Test_INV
xTest_INV5 VDD VSS net4 net5 Test_INV
xTest_INV6 VDD VSS net5 net6 Test_INV
xTest_INV7 VDD VSS net6 OUT Test_INV
**** begin user architecture code

.include /home/shahidosic/OSPDKs/GF180/PDK/share/pdk/gf180mcuC/libs.tech/ngspice/design.spice
.lib /home/shahidosic/OSPDKs/GF180/PDK/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.spice typical



.ic v(OUT)=0
.control
save all
tran 10p 100n
plot v(OUT)
write inv_tb.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/Test_INV.sym # of pins=4
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/Test_INV.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/Test_INV.sch
.subckt Test_INV VDD VSS IN OUT
*.ipin IN
*.iopin VDD
*.iopin VSS
*.opin OUT
XM1 OUT IN VSS VSS nmos_3p3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
