** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/inv_dc_tb.sch
**.subckt inv_dc_tb
C1 OUT VSS 20f m=1
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3
.save i(v2)
V3 IN VSS 3
.save i(v3)
xTest_INV1 VDD VSS IN OUT Test_INV
**** begin user architecture code

.include ./ngspice/design.spice
.lib ./ngspice/sm141064.spice typical



.control
save all
dc V3 0 3 0.01
plot v(IN) v(OUT)
op
write inv_dc_tb.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/Test_INV.sym # of pins=4
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/Test_INV.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/Test_INV.sch
.subckt Test_INV VDD VSS IN OUT
*.ipin IN
*.iopin VDD
*.iopin VSS
*.opin OUT
XM1 OUT IN VSS VSS nmos_3p3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pmos_3p3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
