** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/PLL_COMPLETE.sch
**.subckt PLL_COMPLETE
xPFD1 VDD VSS IN OSCOUTBY64 QA QB PFD
xCP1 VDD IIN5U VBIAS VCTRL IOUT5U VSS RSTB QB QA CP
xVCO1 VDD VSS VBIAS VCTRL net1 VCO
xinv_one1 VDD VSS net1 net2 INV_one
xinv_four1 VDD VSS net2 OSCOUT INV_four
C3 OSCOUT VSS 10f m=1
xFBY641 VDD VSS OSCOUT RSTB OSCOUTBY64 FBY64
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
V3 IN VSS pulse(0 3.3 0 100p 100p 250n 500n)
.save i(v3)
V4 RSTB VSS pwl(0 0 50n 0 51n 3.3 )
.save i(v4)
xBiasGen1 VDD VSS IOUT5U IIN5U IBIAS100U BiasGen
I1 VDD IBIAS100U 100u
xFBY161 VDD VSS OSCOUT VDD net3 FBY16
xFBY321 VDD VSS VDD OSCOUT net4 FBY32
R1 net6 OUTBY16 100 m=1
C1 OUTBY16 VSS 5p m=1
xPAD_DRIVER1 VDD VSS net3 net6 PAD_DRIVER
xPAD_DRIVER2 VDD VSS net4 net5 PAD_DRIVER
R2 net5 OUTBY32 100 m=1
C2 OUTBY32 VSS 5p m=1
**** begin user architecture code

.include /home/shahidosic/OSPDKs/GF180/PDK/share/pdk/gf180mcuC/libs.tech/ngspice/design.spice
.lib /home/shahidosic/OSPDKs/GF180/PDK/share/pdk/gf180mcuC/libs.tech/ngspice/sm141064.spice typical



.ic v(out)=0
.option TEMP=27 wnflag=1
.control
*save all
save v(VCTRL) v(OSCOUT) v(OSCOUTBY64) v(IN) v(QA) v(QB) v(OUTBY16) v(OUTBY32)
tran 20p 50u
*plot v(OUTBY64) v(IN)
plot v(VCTRL) v(OSCOUT)
WRDATA PLL_Complete.csv v(VCTRL) v(OSCOUT) v(OSCOUTBY64) v(IN) v(QA) v(QB) v(OUTBY16) v(OUTBY32)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/PFD.sym # of pins=6
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/PFD.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/PFD.sch
.subckt PFD VDD VSS A B QA QB
*.ipin A
*.iopin VDD
*.iopin VSS
*.opin QA
*.ipin B
*.opin QB
xDFF1 VDD VSS VDD A QA net2 net1 DFF
xDFF2 VDD VSS VDD B QB net3 net1 DFF
xNAND1 VDD VSS QA net1 QB NAND
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/CP.sym # of pins=9
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/CP.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/CP.sch
.subckt CP VDD IIN5U VBIAS VCTRL IOUT5U VSS RSTB QB QA
*.iopin VDD
*.iopin VCTRL
*.ipin RSTB
*.ipin QA
*.ipin QB
*.iopin IIN5U
*.iopin IOUT5U
*.iopin VSS
*.iopin VBIAS
XM1 VBIAS VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM2 VBIAS VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
C2 VBIAS VSS 1p m=1
xinv_one2 VDD VSS QA net2 INV_one
XM3 net3 IOUT5U VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM4 net4 net2 net3 VDD pmos_3p3 L=0.28u W=3u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM5 net4 net1 net5 VSS nmos_3p3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM6 net5 IIN5U VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM7 IOUT5U IOUT5U VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM8 IIN5U IIN5U VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
R1 VCTRL net6 100k m=1
C1 net6 VSS 10p m=1
XM9 net7 RSTB VDD VDD pmos_3p3 L=0.6u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM10 VCTRL RSTB net7 VDD pmos_3p3 L=0.6u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
xTG1 VDD VSS VDD QB net1 TG
xTG2 VDD VSS RSTB net4 VCTRL TG
C4 VCTRL VSS 2p m=1
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/VCO.sym # of pins=5
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/VCO.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/VCO.sch
.subckt VCO VDD VSS VBIAS VCTRL OSC
*.iopin VDD
*.iopin VSS
*.iopin OSC
*.iopin VBIAS
*.iopin VCTRL
XM5 net7 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM3 net8 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM4 net9 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM8 net10 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM9 net11 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM10 net12 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM11 net13 VBIAS VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM6 net14 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM7 net15 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM12 net16 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM13 net17 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM15 net18 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM16 net19 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM17 net20 VCTRL VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
xinv1 net7 net14 OSC net1 inv
xinv2 net8 net15 net1 net2 inv
xinv3 net9 net16 net2 net3 inv
xinv4 net10 net17 net3 net4 inv
xinv5 net11 net18 net4 net5 inv
xinv6 net12 net19 net5 net6 inv
xinv7 net13 net20 net6 OSC inv
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/INV_one.sym # of pins=4
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/INV_one.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/INV_one.sch
.subckt INV_one VDD VSS IN OUT
*.ipin IN
*.iopin VDD
*.iopin VSS
*.opin OUT
XM1 OUT IN VSS VSS nmos_3p3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT IN VDD VDD pmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/INV_four.sym # of pins=4
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/INV_four.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/INV_four.sch
.subckt INV_four VDD VSS IN OUT
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
xinv_one1 VDD VSS IN OUT INV_one
xinv_one2 VDD VSS IN OUT INV_one
xinv_one3 VDD VSS IN OUT INV_one
xinv_one4 VDD VSS IN OUT INV_one
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/FBY64.sym # of pins=5
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/FBY64.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/FBY64.sch
.subckt FBY64 VDD VSS IN RSTB OUT
*.ipin IN
*.iopin VDD
*.iopin VSS
*.opin OUT
*.ipin RSTB
xDFF1 VDD VSS net1 IN net2 net1 RSTB DFF
xDFF2 VDD VSS net3 net2 net4 net3 RSTB DFF
xDFF3 VDD VSS net5 net4 net6 net5 RSTB DFF
xDFF4 VDD VSS net7 net6 net8 net7 RSTB DFF
xDFF5 VDD VSS net9 net8 net10 net9 RSTB DFF
xDFF6 VDD VSS net11 net10 OUT net11 RSTB DFF
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/BiasGen.sym # of pins=5
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/BiasGen.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/BiasGen.sch
.subckt BiasGen VDD VSS IOUT5U IIN5U IBIAS100U
*.iopin VDD
*.iopin IIN5U
*.iopin IOUT5U
*.iopin VSS
*.iopin IBIAS100U
XM7 net2 net2 VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM8 VB VB VSS VSS nmos_3p3 L=0.6u W=100u nf=20 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM1 net1 VB VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 net5 net2 VDD VDD pmos_3p3 L=0.6u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net3 VB VSS VSS nmos_3p3 L=0.6u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 IBIAS100U IBIAS100U VB VSS nmos_3p3 L=0.6u W=125u nf=25 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 net4 IBIAS100U net1 VSS nmos_3p3 L=0.6u W=10u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net4 net4 net2 VDD pmos_3p3 L=0.6u W=30u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM9 IIN5U net4 net5 VDD pmos_3p3 L=0.6u W=30u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM10 IOUT5U IBIAS100U net3 VSS nmos_3p3 L=0.6u W=10u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/FBY16.sym # of pins=5
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/FBY16.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/FBY16.sch
.subckt FBY16 VDD VSS IN RSTB OUT
*.ipin IN
*.iopin VDD
*.iopin VSS
*.opin OUT
*.ipin RSTB
xDFF1 VDD VSS net1 IN net2 net1 RSTB DFF
xDFF2 VDD VSS net3 net2 net4 net3 RSTB DFF
xDFF3 VDD VSS net5 net4 net6 net5 RSTB DFF
xDFF4 VDD VSS net7 net6 OUT net7 RSTB DFF
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/FBY32.sym # of pins=5
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/FBY32.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/FBY32.sch
.subckt FBY32 VDD VSS IN RSTB OUT
*.ipin IN
*.iopin VDD
*.iopin VSS
*.opin OUT
*.ipin RSTB
xDFF1 VDD VSS net1 IN net2 net1 RSTB DFF
xDFF2 VDD VSS net3 net2 net4 net3 RSTB DFF
xDFF3 VDD VSS net5 net4 net6 net5 RSTB DFF
xDFF4 VDD VSS net7 net6 net8 net7 RSTB DFF
xDFF5 VDD VSS net9 net8 OUT net9 RSTB DFF
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/PAD_DRIVER.sym # of pins=4
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/PAD_DRIVER.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/PAD_DRIVER.sch
.subckt PAD_DRIVER VDD VSS IN OUT
*.iopin VDD
*.opin OUT
*.ipin IN
*.iopin VSS
xinv_four1 VDD VSS IN net1 INV_four
xinv_sixteen1 VDD VSS net1 OUT INV_sixteen
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/DFF.sym # of pins=7
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/DFF.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/DFF.sch
.subckt DFF VDD VSS D CLK Q QB RSTB
*.ipin D
*.iopin VDD
*.iopin VSS
*.opin Q
*.ipin CLK
*.opin QB
*.ipin RSTB
xNAND2 VDD VSS net1 net4 net3 NAND
xNAND_TI1 VDD VSS net4 net3 RSTB CLK NAND_TI
xNAND_TI2 VDD VSS net3 net2 net1 CLK NAND_TI
xNAND_TI3 VDD VSS net2 net1 D RSTB NAND_TI
xNAND3 VDD VSS net3 Q QB NAND
xNAND_TI4 VDD VSS Q QB net2 RSTB NAND_TI
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/NAND.sym # of pins=5
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/NAND.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/NAND.sch
.subckt NAND VDD VSS A OUT B
*.ipin A
*.iopin VDD
*.iopin VSS
*.opin OUT
*.ipin B
XM1 OUT A net1 VSS nmos_3p3 L=0.28u W=1.6u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT A VDD VDD pmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 B VSS VSS nmos_3p3 L=0.28u W=1.6u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 OUT B VDD VDD pmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/TG.sym # of pins=5
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/TG.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/TG.sch
.subckt TG VDD VSS CLK A B
*.iopin A
*.iopin VDD
*.iopin VSS
*.iopin B
*.ipin CLK
XM3 A CLKB B VDD pmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 A CLK B VSS nmos_3p3 L=0.28u W=0.8u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
xinv_one1 VDD VSS CLK CLKB INV_one
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/inv.sym # of pins=4
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/inv.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/inv.sch
.subckt inv VDD VSS IN OUT
*.ipin IN
*.iopin VDD
*.iopin VSS
*.opin OUT
XM1 OUT IN VSS VSS nmos_3p3 L=1u W=5u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
XM2 OUT IN VDD VDD pmos_3p3 L=1u W=15u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=2
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/INV_sixteen.sym # of pins=4
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/INV_sixteen.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/INV_sixteen.sch
.subckt INV_sixteen VDD VSS IN OUT
*.iopin VDD
*.iopin VSS
*.ipin IN
*.opin OUT
xinv_four1 VDD VSS IN OUT INV_four
xinv_four2 VDD VSS IN OUT INV_four
xinv_four3 VDD VSS IN OUT INV_four
xinv_four4 VDD VSS IN OUT INV_four
.ends


* expanding   symbol:  /home/shahidosic/GFProjects/PLL/Xschem/NAND_TI.sym # of pins=6
** sym_path: /home/shahidosic/GFProjects/PLL/Xschem/NAND_TI.sym
** sch_path: /home/shahidosic/GFProjects/PLL/Xschem/NAND_TI.sch
.subckt NAND_TI VDD VSS A OUT C B
*.ipin A
*.iopin VDD
*.iopin VSS
*.opin OUT
*.ipin B
*.ipin C
XM1 OUT A net1 VSS nmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM2 OUT A VDD VDD pmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM3 net1 B net2 VSS nmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM4 OUT B VDD VDD pmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM5 OUT C VDD VDD pmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
XM6 net2 C VSS VSS nmos_3p3 L=0.28u W=2.4u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
